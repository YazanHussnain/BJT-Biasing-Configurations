FIXED BIAS CONFIGURATION
*Title Line
VCC 1 0 15
*15V Voltage source
RC 1 3 7.5k
RB 1 2 1430k
.model 2N3904 NPN(Is=6.734f Xti=3 Eg=1.11 Vaf=74.03 Bf=416.4 Ne=1.259
+               Ise=6.734f Ikf=66.78m Xtb=1.5 Br=.7371 Nc=2 Isc=0 Ikr=0 Rc=1
+               Cjc=3.638p Mjc=.3085 Vjc=.75 Fc=.5 Cje=4.493p Mje=.2593 Vje=.75
+               Tr=239.5n Tf=301.2p Itf=.4 Vtf=4 Xtf=2 Rb=10)
Q1 3 2 0 2N3904
* Connect BJT at nodes 3, 2, 0
.TRAN 1NS 700NS 0NS
* Transient Analysis
.PLOT TRAN V(3,0)
* Plot graph of V(3) - V(0)
.OP
* Give voltage at each and node and current in each branch
.END